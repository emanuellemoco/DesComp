library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;           

entity projeto1 is
    port(
        SW: in std_logic_vector(9 downto 0);
        LEDR: out std_logic_vector(9 downto 0);
        KEY: in std_logic_vector(3 downto 0);
		CLOCK_50: in std_logic;
		FPGA_RESET_n: in std_logic
);
end entity;

architecture arch of projeto1 is

    component registradorGenerico is
        generic (
            larguraDados : natural := 8
        );
        port (DIN : in std_logic_vector(larguraDados-1 downto 0);
           DOUT : out std_logic_vector(larguraDados-1 downto 0);
           ENABLE : in std_logic;
           CLK,RST : in std_logic
            );
    end component;

    component mux2x1 is
        generic (
			larguraDados : natural := 8
		);
        port (
            entradaA_MUX, entradaB_MUX : in std_logic_vector((larguraDados-1) downto 0);
            seletor_MUX : in std_logic;
            saida_MUX : out std_logic_vector((larguraDados-1) downto 0)
          );
    end component; 

    component ULAsoma is
        generic ( larguraDados : natural := 8);
        port (
          entradaA, entradaB: in STD_LOGIC_VECTOR((larguraDados-1) downto 0);
          operacao: in STD_LOGIC;
          saida: out STD_LOGIC_VECTOR((larguraDados-1) downto 0)
        );
      end component;



    component edgeDetector is
        Port ( clk     : in  STD_LOGIC;
                 entrada : in  STD_LOGIC;
                 saida   : out STD_LOGIC);
   end component;

SIGNAL muxOut, regAout, regBout, ulaOut: std_logic_vector( 7 downto 0); 
SIGNAL rstAOut, rstBOut, clkOut: std_logic;

begin

    detectorCLK: edgeDetector  port map (CLOCK_50, FPGA_RESET_N, clkOut);

    detectorRSTA: edgeDetector  port map (CLOCK_50, KEY(1), rstAOut);

    detectorRSTB: edgeDetector  port map (CLOCK_50, KEY(0), rstBOut);

    muxIN_A: mux2x1 port map (SW(7 downto 0), ulaOut, SW(8), muxOut);

    regA: registradorGenerico port map (muxOut, regAout, KEY(3), clkOut, rstAOut);

    regB: registradorGenerico port map (SW(7 downto 0), regBout, KEY(2), clkOut, rstBOut);

    ULA: ULAsoma port map (regAOut, regBOut, SW(9), ulaOut);

	LEDR <= SW(9 downto 8) & ulaOut ;
		  
end architecture;